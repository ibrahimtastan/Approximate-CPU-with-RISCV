`timescale 100ps / 1ps

module buffer_cell(
	input in1,in2,
	output out1,out2
    );

assign out1 = in1;
assign out2 = in2;

endmodule
